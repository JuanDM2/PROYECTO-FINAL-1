library verilog;
use verilog.vl_types.all;
entity Output_ports_vlg_vec_tst is
end Output_ports_vlg_vec_tst;
